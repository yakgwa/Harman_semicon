`timescale 1ns / 1ps

module ROM (
    input  logic [31:0] addr,
    output logic [31:0] data
);
    logic [31:0] rom[0:2**8-1];

    initial begin
        //$readmemh("code_mem1.mem", rom);
        // R - funct7, rs2, rs1, funct3, rd, opcode
        rom[0] = 32'b0000000_00001_00010_000_00100_0110011; // add x4, x2, x1
        rom[1] = 32'b0100000_00001_00010_000_00101_0110011; // sub x5, x2, x1
        rom[2] = 32'b0000000_00000_00011_111_00110_0110011; // and x6, x3, x0
        rom[3] = 32'b0000000_00000_00011_110_00111_0110011; // or x7, x3, x0
        // I - imm, rs1, funct3, rd, opcode
        rom[4] = 32'b000000000001_00001_000_01001_0010011; // addi x9, x1, 1
        rom[5] = 32'b000000000100_00010_111_01010_0010011; // andi x10, x2, 4
        rom[6] = 32'b000000000011_00001_001_01011_0010011; // slli x11, x1, 3
        // S - imm7, rs2, rs1, funct3, imm5, opcode
        rom[7] = 32'b0000000_00001_01100_000_00000_0100011; // sb x1, x12, 0
        rom[8] = 32'b0000000_00001_01101_001_00000_0100011; // sh x1, x13, 0
        rom[9] = 32'b0000000_00001_01110_010_00000_0100011; // sw x1, x14, 0
        //rom[10] = 32'b0000000_00010_01111_010_00000_0100011; // sw x3, x15, 0
        //rom[11] = 32'b0000000_00010_01111_010_00011_0100011; // sw x2, x15, 3
        // B - imm7, rs2, rs1, funct3, imm5, opcode
        rom[10] = 32'b0000000_00010_00010_000_01000_1100011; // beq x2, x2, 8 (2 Shift)
        rom[12] = 32'b0000000_00010_00011_001_01100_1100011; // bne x2, x3, 12  
        //rom[12] = 32'b0000000_00010_00010_000_00100_1100011; // blt x2, x2, 12      
        // L - imm12, rs1, funct3, rs2, opcode
        rom[13] = 32'b000000000000_01110_000_10000_0000011; // lb x16, 0(x14)
        rom[14] = 32'b000000000000_01110_001_10001_0000011; // lh x17, 0(x14)
        rom[15] = 32'b000000000000_01110_010_10010_0000011; // lw x18, 0(x14)
        rom[16] = 32'b000000000000_01110_100_10011_0000011; // lbu x19, 0(x14)
        rom[17] = 32'b000000000000_01110_101_10100_0000011; // lhu x20, 0(x14)
        // LU - imm20, rd, opcode
        rom[18] = 32'b00010000000000000000_10101_0110111; // lui x21, x10000000;
        // AU - imm20, rd, opcode
        rom[19] = 32'b10101011110011011110_10110_0010111; //auipc 0xABCDE (Plus 12 & Store x22)
        // J - imm20, rd, opcode
        // rom[20] = 32'b1_1111111100_1_11111111_00000_1101111; // jal x0, -8;        
        // JL - imm20, rs1, funct3, rd, opcode
        rom[20] = 32'b000000000100_00010_000_10111_1100111; // jarl x23, x2, 8 (rd : x23, jump addr = x2 + 4)

    end

    assign data = rom[addr[31:2]];
endmodule
