`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/10/13 14:39:00
// Design Name: 
// Module Name: tb_rv32i
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_rv32i();
    logic clk;
    logic reset;

    MCU dut(.*);

    always #5 clk = ~clk;

    initial begin
        #00 clk = 0; reset = 1;
        #10 reset = 0;
        #3000 $finish;
    end

endmodule
