`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/09/02 17:54:50
// Design Name: 
// Module Name: button_debounce_ori
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module button_debounce_ori(
    input clk, rst,
    input i_btn,
    output o_btn
    );

    // 100m -> 1m
    reg[$clog2(100)-1:0] counter_reg;
    reg clk_reg;
    reg [7:0] q_reg, q_next;
    reg edge_reg;
    wire debounce;

    // clock divider
    always@(posedge clk or posedge rst) begin
        if(rst) begin
            counter_reg <= 0;
            clk_reg <= 1'b0;
        end else begin
            if(counter_reg == 99) begin
                counter_reg <= 0;
                clk_reg <= 1'b1;
            end else begin
                counter_reg <= counter_reg + 1;
                clk_reg <= 1'b0;
            end
        end
    end

    // debounce logic, shift register
    always @(posedge clk_reg or posedge rst) begin
        if(rst) begin
            q_reg <= 0;//4'b0;
        end else begin
            q_reg <= q_next; 
        end    
    end

    // Serial input, Paraller output shift register
    always@(*) begin
        q_next = {i_btn, q_reg[7:1]}; //q_reg[3:1]};
   
    end

    assign debounce = &q_reg; 

    // Q5 output
    always@(posedge clk or posedge rst) begin
        if(rst) begin
            edge_reg <= 1'b0;
        end else begin
            edge_reg <= debounce;
        end
    end

    // edge output
    assign o_btn = ~edge_reg & debounce;


endmodule
